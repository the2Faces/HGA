LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY HGA IS

PORT
(
	KMM, KOM, MIL, E_STOP : IN STD_LOGIC;
	KAV, MIV : OUT STD_LOGIC;
	clk : IN STD_LOGIC;
	START , out_50_50 : OUT STD_LOGIC;
	A_STOP, POR : IN STD_LOGIC
);

END ENTITY HGA;

ARCHITECTURE beh OF HGA IS

TYPE states IS (IGZ );
SIGNAL current_state, next_state : states;



BEGIN



END ARCHITECTURE beh;