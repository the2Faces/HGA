LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY LTVC IS
PORT
(
	KAV, MIV : IN STD_LOGIC;
	KON, MON : OUT STD_LOGIC
);
END ENTITY LTVC;

ARCHITECTURE beh OF LTVC is
BEGIN

KON <= KAV;
MON <= MIV;

END ARCHITECTURE beh;