LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY HGA IS

PORT
(
	KMM, KOM, MIL, E_STOP : IN STD_LOGIC;
	A_STOP, POR : OUT STD_LOGIC
);

END ENTITY HGA;

ARCHITECTURE beh OF HGA IS

SIGNAL test2sig : STD_LOGIC;
SIGNAL inttest : STD_LOGIC;
BEGIN



END ARCHITECUTRE beh OF HGA;